CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
21
10 3-In NAND~
219 882 605 0 4 22
0 3 4 5 7
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U8A
263 -528 284 -520
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 8 0
1 U
5130 0 0
2
5.89972e-315 5.32571e-315
0
10 3-In NAND~
219 883 672 0 4 22
0 5 4 2 6
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U4C
-15 -183 6 -175
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 4 0
1 U
391 0 0
2
5.89972e-315 5.30499e-315
0
10 2-In NAND~
219 1058 687 0 3 22
0 3 6 2
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7B
71 -589 92 -581
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3124 0 0
2
5.89972e-315 5.26354e-315
0
10 2-In NAND~
219 1055 589 0 3 22
0 7 2 3
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7A
37 -461 58 -453
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3421 0 0
2
5.89972e-315 0
0
10 3-In NAND~
219 797 282 0 4 22
0 11 10 8 14
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U4A
323 -249 344 -241
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
8157 0 0
2
5.89972e-315 5.32571e-315
0
10 3-In NAND~
219 798 349 0 4 22
0 8 9 12 13
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U4B
341 -272 362 -264
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 4 0
1 U
5572 0 0
2
5.89972e-315 5.30499e-315
0
10 2-In NAND~
219 973 364 0 3 22
0 12 13 11
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3C
177 -279 198 -271
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8901 0 0
2
5.89972e-315 5.26354e-315
0
10 2-In NAND~
219 970 266 0 3 22
0 14 11 12
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3D
177 -211 198 -203
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7361 0 0
2
5.89972e-315 0
0
9 Inverter~
13 190 638 0 2 22
0 15 16
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U6A
921 -586 942 -578
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
4747 0 0
2
5.89972e-315 0
0
10 2-In NAND~
219 318 611 0 3 22
0 15 17 21
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5D
-163 -131 -142 -123
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
972 0 0
2
5.89972e-315 5.32571e-315
0
10 2-In NAND~
219 319 663 0 3 22
0 17 16 20
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5C
-127 -179 -106 -171
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3472 0 0
2
5.89972e-315 5.30499e-315
0
10 2-In NAND~
219 490 599 0 3 22
0 21 18 19
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5B
-239 -94 -218 -86
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9998 0 0
2
5.89972e-315 5.26354e-315
0
10 2-In NAND~
219 494 672 0 3 22
0 19 20 18
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5A
-313 -180 -292 -172
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3536 0 0
2
5.89972e-315 0
0
10 2-In NAND~
219 495 451 0 3 22
0 23 27 22
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4597 0 0
2
5.89972e-315 0
0
10 2-In NAND~
219 492 353 0 3 22
0 28 22 23
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3835 0 0
2
5.89972e-315 0
0
10 2-In NAND~
219 322 436 0 3 22
0 24 25 27
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3670 0 0
2
5.89972e-315 0
0
10 2-In NAND~
219 318 369 0 3 22
0 26 24 28
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5616 0 0
2
5.89972e-315 0
0
9 2-In NOR~
219 659 184 0 3 22
0 29 31 30
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9323 0 0
2
5.89972e-315 0
0
9 2-In NOR~
219 657 110 0 3 22
0 32 30 29
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
317 0 0
2
5.89972e-315 0
0
10 2-In NAND~
219 205 192 0 3 22
0 34 35 33
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3108 0 0
2
5.89972e-315 0
0
10 2-In NAND~
219 202 104 0 3 22
0 36 33 34
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4299 0 0
2
5.89972e-315 0
0
51
0 3 2 0 0 8320 0 0 2 9 0 5
1096 687
1096 707
829 707
829 681
859 681
0 1 3 0 0 8320 0 0 1 10 0 5
1092 589
1092 568
821 568
821 596
858 596
0 2 4 0 0 4096 0 0 2 5 0 3
816 605
816 672
859 672
0 2 5 0 0 4224 0 0 0 0 6 2
777 638
851 638
0 2 4 0 0 4224 0 0 1 0 0 2
787 605
858 605
3 1 5 0 0 0 0 1 2 0 0 4
858 614
851 614
851 663
859 663
2 0 2 0 0 0 0 4 0 0 9 5
1031 598
996 598
996 642
1103 642
1103 687
0 1 3 0 0 0 0 0 3 10 0 5
1103 589
1103 624
985 624
985 678
1034 678
3 2 2 0 0 0 0 3 0 0 0 2
1085 687
1161 687
2 3 3 0 0 0 0 0 4 0 0 2
1154 589
1082 589
4 2 6 0 0 12416 0 2 3 0 0 4
910 672
964 672
964 696
1034 696
4 1 7 0 0 12416 0 1 4 0 0 4
909 605
964 605
964 580
1031 580
0 2 8 0 0 4224 0 0 0 0 18 2
692 315
766 315
0 2 9 0 0 4224 0 0 6 0 0 2
699 349
774 349
0 2 10 0 0 4224 0 0 5 0 0 2
702 282
773 282
0 1 11 0 0 8320 0 0 5 21 0 5
1049 364
1049 244
738 244
738 273
773 273
0 3 12 0 0 8320 0 0 6 22 0 5
1038 266
1038 384
738 384
738 358
774 358
3 1 8 0 0 0 0 5 6 0 0 4
773 291
766 291
766 340
774 340
2 0 11 0 0 0 0 8 0 0 21 5
946 275
911 275
911 319
1018 319
1018 364
0 1 12 0 0 0 0 0 7 22 0 5
1018 266
1018 301
900 301
900 355
949 355
3 2 11 0 0 0 0 7 0 0 0 2
1000 364
1076 364
2 3 12 0 0 0 0 0 8 0 0 2
1069 266
997 266
4 2 13 0 0 12416 0 6 7 0 0 4
825 349
879 349
879 373
949 373
4 1 14 0 0 12416 0 5 8 0 0 4
824 282
879 282
879 257
946 257
0 2 15 0 0 4096 0 0 0 0 27 2
147 601
193 601
2 2 16 0 0 8320 0 9 11 0 0 3
193 656
193 672
295 672
1 1 15 0 0 4224 0 10 9 0 0 5
294 602
193 602
193 595
193 595
193 620
0 2 17 0 0 4224 0 0 0 0 35 2
235 639
280 639
2 0 18 0 0 12416 0 12 0 0 31 5
466 608
432 608
432 641
539 641
539 673
0 1 19 0 0 8320 0 0 13 32 0 5
539 599
539 623
421 623
421 663
470 663
3 2 18 0 0 0 0 13 0 0 0 4
521 672
539 672
539 673
597 673
2 3 19 0 0 0 0 0 12 0 0 2
590 599
517 599
3 2 20 0 0 12416 0 11 13 0 0 4
346 663
400 663
400 681
470 681
3 1 21 0 0 12416 0 10 12 0 0 4
345 611
400 611
400 590
466 590
2 1 17 0 0 0 0 10 11 0 0 4
294 620
280 620
280 654
295 654
2 0 22 0 0 12416 0 15 0 0 38 5
468 362
433 362
433 406
540 406
540 451
0 1 23 0 0 8320 0 0 14 39 0 5
540 353
540 388
422 388
422 442
471 442
3 2 22 0 0 0 0 14 0 0 0 2
522 451
598 451
2 3 23 0 0 0 0 0 15 0 0 2
591 353
519 353
0 1 26 0 0 4224 0 0 17 0 0 2
221 360
294 360
3 2 27 0 0 12416 0 16 14 0 0 4
349 436
401 436
401 460
471 460
3 1 28 0 0 12416 0 17 15 0 0 4
345 369
401 369
401 344
468 344
2 1 24 0 0 0 0 17 16 0 0 4
294 378
285 378
285 427
298 427
1 0 29 0 0 12416 0 18 0 0 47 5
646 175
601 175
601 140
719 140
719 110
2 0 30 0 0 12416 0 19 0 0 46 5
644 119
582 119
582 154
722 154
722 184
3 2 30 0 0 0 0 18 0 0 0 2
698 184
771 184
3 2 29 0 0 0 0 19 0 0 0 2
696 110
771 110
2 0 33 0 0 12288 0 21 0 0 50 5
178 113
148 113
148 152
268 152
268 192
0 1 34 0 0 8192 0 0 20 51 0 5
269 104
269 132
160 132
160 183
181 183
3 0 33 0 0 4224 0 20 0 0 0 3
232 192
384 192
384 185
3 0 34 0 0 4224 0 21 0 0 0 3
229 104
383 104
383 100
35
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
581 315 610 339
591 323 599 339
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
586 419 615 443
596 427 604 443
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
581 337 610 361
591 345 599 361
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
587 436 616 460
597 444 605 460
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
582 406 619 430
592 414 608 430
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
583 629 620 653
593 637 609 653
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
586 658 615 682
596 666 604 682
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
579 582 608 606
589 590 597 606
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
586 643 615 667
596 651 604 667
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
581 596 610 620
591 604 599 620
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
223 624 252 648
233 632 241 648
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
197 623 242 647
207 631 231 647
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
134 586 163 610
144 594 152 610
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
137 572 162 596
145 580 153 596
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
681 299 710 323
691 307 699 323
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
654 302 699 326
664 310 688 326
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
667 334 696 358
677 342 685 358
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
683 333 712 357
693 341 701 357
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
666 265 695 289
676 273 684 289
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
684 266 713 290
694 274 702 290
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1059 228 1088 252
1069 236 1077 252
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1064 332 1093 356
1074 340 1082 356
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1059 250 1088 274
1069 258 1077 274
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1065 349 1094 373
1075 357 1083 373
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1060 319 1097 343
1070 327 1086 343
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
766 622 795 646
776 630 784 646
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
739 625 784 649
749 633 773 649
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
569 696 598 720
579 704 587 720
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1144 551 1173 575
1154 559 1162 575
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1149 655 1178 679
1159 663 1167 679
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1144 573 1173 597
1154 581 1162 597
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1150 672 1179 696
1160 680 1168 696
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1145 642 1182 666
1155 650 1171 666
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
769 589 794 613
777 597 785 613
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
751 588 776 612
759 596 767 612
1 T
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
