CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 580 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
22
14 Logic Display~
6 594 898 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
44395.7 0
0
9 2-In AND~
219 326 891 0 3 22
0 9 8 13
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3670 0 0
2
44395.7 7
0
9 2-In AND~
219 367 954 0 3 22
0 10 11 12
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5616 0 0
2
44395.7 6
0
9 2-In XOR~
219 268 963 0 3 22
0 9 8 11
0
0 0 608 0
5 74F86
-18 -24 17 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9323 0 0
2
44395.7 5
0
8 2-In OR~
219 476 920 0 3 22
0 13 12 7
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
317 0 0
2
44395.7 4
0
13 Logic Switch~
5 135 854 0 1 11
0 10
0
0 0 21344 0
2 0V
-32 -5 -18 3
2 V9
1030 510 1044 518
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3108 0 0
2
44395.7 2
0
13 Logic Switch~
5 136 882 0 1 11
0 8
0
0 0 21344 0
2 0V
-30 -5 -16 3
2 V8
1034 471 1048 479
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4299 0 0
2
44395.7 1
0
13 Logic Switch~
5 135 915 0 1 11
0 9
0
0 0 21344 0
2 0V
-30 -4 -16 4
2 V7
1037 431 1051 439
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9672 0 0
2
44395.7 0
0
13 Logic Switch~
5 142 531 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-32 -5 -18 3
2 V6
1030 510 1044 518
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7876 0 0
2
44395.7 0
0
13 Logic Switch~
5 143 559 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-30 -5 -16 3
2 V5
1034 471 1048 479
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6369 0 0
2
44395.7 1
0
13 Logic Switch~
5 142 592 0 1 11
0 6
0
0 0 21344 0
2 0V
-30 -4 -16 4
2 V4
1037 431 1051 439
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9172 0 0
2
44395.7 2
0
13 Logic Switch~
5 100 165 0 1 11
0 9
0
0 0 21344 0
2 0V
-30 -4 -16 4
2 V3
1037 431 1051 439
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7100 0 0
2
44395.7 3
0
13 Logic Switch~
5 101 132 0 1 11
0 8
0
0 0 21344 0
2 0V
-30 -5 -16 3
2 V2
1034 471 1048 479
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3820 0 0
2
44395.7 4
0
13 Logic Switch~
5 100 104 0 1 11
0 10
0
0 0 21344 0
2 0V
-32 -5 -18 3
2 V1
1030 510 1044 518
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7678 0 0
2
44395.7 5
0
8 2-In OR~
219 491 627 0 3 22
0 6 3 2
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
961 0 0
2
44395.7 6
0
14 Logic Display~
6 604 623 0 1 2
10 2
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
44395.7 7
0
9 2-In NOR~
219 313 659 0 3 22
0 5 4 3
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3409 0 0
2
44395.7 8
0
14 Logic Display~
6 757 286 0 1 2
10 7
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
44395.7 9
0
8 2-In OR~
219 604 290 0 3 22
0 13 12 7
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8885 0 0
2
44395.7 10
0
9 2-In XOR~
219 310 358 0 3 22
0 9 8 11
0
0 0 608 0
5 74F86
-18 -24 17 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3780 0 0
2
44395.7 11
0
9 2-In AND~
219 452 336 0 3 22
0 10 11 12
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9265 0 0
2
44395.7 12
0
9 2-In AND~
219 383 240 0 3 22
0 9 8 13
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9442 0 0
2
44395.7 13
0
23
3 1 0 0 0 0 0 5 1 0 0 3
509 920
594 920
594 916
3 2 0 0 0 0 0 3 5 0 0 4
388 954
410 954
410 929
463 929
1 1 0 0 0 0 0 6 3 0 0 6
147 854
164 854
164 923
310 923
310 945
343 945
3 2 0 0 0 0 0 4 3 0 0 2
301 963
343 963
3 1 0 0 0 0 0 2 5 0 0 4
347 891
398 891
398 911
463 911
0 2 0 0 0 0 0 0 4 8 0 3
184 882
184 972
252 972
0 1 0 0 0 0 0 0 4 9 0 3
200 915
200 954
252 954
1 1 0 0 0 0 0 7 2 0 0 2
148 882
302 882
1 2 0 0 0 0 0 8 2 0 0 4
147 915
222 915
222 900
302 900
3 1 2 0 0 4224 0 15 16 0 0 2
524 627
588 627
3 2 3 0 0 12416 0 17 15 0 0 4
352 659
410 659
410 636
478 636
1 2 4 0 0 8320 0 9 17 0 0 4
154 531
194 531
194 668
300 668
1 1 5 0 0 12416 0 10 17 0 0 4
155 559
175 559
175 650
300 650
1 1 6 0 0 8320 0 11 15 0 0 3
154 592
154 618
478 618
1 3 7 0 0 4224 0 18 19 0 0 2
741 290
637 290
2 0 8 0 0 4096 0 22 0 0 19 2
359 249
131 249
1 0 9 0 0 4224 0 22 0 0 20 2
359 231
112 231
1 1 10 0 0 12416 0 14 21 0 0 4
112 104
152 104
152 327
428 327
1 2 8 0 0 8320 0 13 20 0 0 4
113 132
131 132
131 367
294 367
1 1 9 0 0 0 0 12 20 0 0 3
112 165
112 349
294 349
2 3 11 0 0 4224 0 21 20 0 0 4
428 345
351 345
351 358
343 358
3 2 12 0 0 4224 0 21 19 0 0 4
473 336
532 336
532 299
591 299
3 1 13 0 0 4224 0 22 19 0 0 4
404 240
533 240
533 281
591 281
64
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
243 855 270 877
252 863 260 879
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
518 894 577 916
527 901 567 917
5 pin-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
414 931 473 953
423 938 463 954
5 Pin-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
404 886 463 908
413 893 453 909
5 Pin-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
338 865 397 887
347 872 387 888
5 pin-3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
252 896 311 918
261 903 301 919
5 Pin-2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
65 899 110 923
75 907 99 923
3 A =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
65 867 110 891
75 875 99 891
3 B =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
64 836 109 860
74 844 98 860
3 C =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
325 569 380 593
332 575 372 591
5 C = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
324 549 379 573
331 555 371 571
5 B = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
618 614 673 638
625 619 665 635
5 Y = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
251 525 380 546
259 532 371 547
14 INPUT    A = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
245 149 302 170
253 156 293 171
5 C = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
245 126 302 147
253 133 293 148
5 B = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
538 612 585 636
545 618 577 634
4 ____
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
353 688 400 712
360 694 392 710
4 ____
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
349 615 396 639
356 621 388 637
4 ____
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
344 632 399 656
351 637 391 653
5 (A+B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
516 629 587 653
523 635 579 651
7 A+(B+C)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
346 659 409 683
353 665 401 681
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
227 623 290 647
234 629 282 645
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
229 664 292 688
236 669 284 685
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
514 600 577 624
521 605 569 621
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
402 592 465 616
409 597 457 613
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
209 702 324 723
218 709 314 724
12 EXPRESSION :
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
197 594 220 615
204 601 212 616
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
170 325 193 346
177 332 185 347
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
195 663 218 684
202 670 210 685
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
153 294 176 315
160 301 168 316
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
195 625 220 646
203 632 211 647
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
171 364 196 385
179 371 187 386
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
403 339 426 360
410 346 418 361
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
615 564 684 588
625 572 673 588
6 OUTPUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
72 576 117 600
82 584 106 600
3 A =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
72 542 117 566
82 550 106 566
3 B =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
71 513 116 537
81 521 105 537
3 C =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
177 102 298 123
185 108 289 123
13 INPUT   A = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
773 275 832 296
782 282 822 297
5 Y = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
767 189 836 213
777 197 825 213
6 OUTPUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
264 405 421 429
274 413 410 429
17 Y = AB+C(A XOR B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
164 404 265 428
174 412 254 428
10 Expression
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
535 312 612 336
545 320 601 336
7 Pin - 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
242 244 319 268
252 252 308 268
7 Pin - 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
530 232 607 256
540 240 596 256
7 Pin - 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
242 204 319 228
252 212 308 228
7 Pin - 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
344 340 373 364
354 348 362 364
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
355 300 432 324
365 308 421 324
7 Pin - 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
206 363 283 387
216 371 272 387
7 Pin - 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
205 325 282 349
215 333 271 349
7 Pin - 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
454 344 555 368
464 352 544 368
10 C(A XOR B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
617 295 758 319
627 303 747 319
15 Y=AB+C(A XOR B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
638 259 715 283
648 267 704 283
7 Pin - 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
461 309 538 333
471 317 527 333
7 Pin - 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
430 213 507 237
440 221 496 237
7 Pin - 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
29 86 74 110
39 94 63 110
3 C =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
30 117 75 141
40 125 64 141
3 B =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
30 149 75 173
40 157 64 173
3 A =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
168 200 197 224
178 208 186 224
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
171 246 200 270
181 254 189 270
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
388 247 425 271
398 255 414 271
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
315 367 392 391
325 375 381 391
7 A XOR B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
316 705 403 729
323 711 395 727
9 Y=A+(B+C)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
410 632 473 656
417 637 465 653
6 Pin- 2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
